#SpecName      geometry     potential well depth     collision diameter     dipole moment     polarizability     rotational relaxation number
AR                 0   136.500     3.330     0.000     0.000     0.000
N2                 1    97.530     3.621     0.000     1.760     4.000
HE                 0    10.200     2.576     0.000     0.000     0.000
H2                 1    38.000     2.920     0.000     0.790   280.000
H                  0   145.000     2.050     0.000     0.000     0.000
O2                 1   107.400     3.458     0.000     1.600     3.800
O                  0    80.000     2.750     0.000     0.000     0.000
H2O                2   572.400     2.605     1.844     0.000     4.000
OH                 1    80.000     2.750     0.000     0.000     0.000
H2O2               2   107.400     3.458     0.000     0.000     3.800
HO2                2   107.400     3.458     0.000     0.000     1.000
CO                 1    98.100     3.650     0.000     1.950     1.800
CO2                1   244.000     3.763     0.000     2.650     2.100
HOCO               2   498.000     3.590     0.000     0.000     2.000
CH4                2   141.400     3.746     0.000     2.600    13.000
CH3                1   144.000     3.800     0.000     0.000     0.000
CH2                1   144.000     3.800     0.000     0.000     0.000
CH2(S)             1   144.000     3.800     0.000     0.000     0.000
C                  0    71.400     3.298     0.000     0.000     0.000
CH                 1    80.000     2.750     0.000     0.000     0.000
CH3O2H             2   481.800     3.626     0.000     0.000     1.000
CH3O2              2   481.800     3.626     0.000     0.000     1.000 
CH3OH              2   481.800     3.626     0.000     0.000     1.000
CH3O               2   417.000     3.690     1.700     0.000     2.000
CH2OH              2   417.000     3.690     1.700     0.000     2.000
CH2O               2   498.000     3.590     0.000     0.000     2.000
HCO                2   498.000     3.590     0.000     0.000     0.000
HO2CHO             2   436.000     3.970     0.000     0.000     2.000
HOCHO              2   436.000     3.970     0.000     0.000     2.000
OCHO               2   498.000     3.590     0.000     0.000     2.000
C2H6               2   247.500     4.350     0.000     0.000     1.500
C2H5               2   247.500     4.350     0.000     0.000     1.500
C2H5O2H            2   470.600     4.410     0.000     0.000     1.500
C2H5O2             2   470.600     4.410     0.000     0.000     1.500
C2H4               2   238.400     3.496     0.000     0.000     1.500
C2H3               2   265.300     3.721     0.000     0.000     1.000
C2H2               1   265.300     3.721     0.000     0.000     2.500
C2H                1   265.300     3.721     0.000     0.000     2.500
C2H5OH             2   470.600     4.410     0.000     0.000     1.500
C2H5O              2   470.600     4.410     0.000     0.000     1.500
PC2H4OH            2   470.600     4.410     0.000     0.000     1.500
SC2H4OH            2   470.600     4.410     0.000     0.000     1.500
C2H4O2H            2   470.600     4.410     0.000     0.000     1.500
C2H4O1-2           2   436.000     3.970     0.000     0.000     2.000
C2H3O1-2           2   436.000     3.970     0.000     0.000     2.000
CH3CHO             2   436.000     3.970     0.000     0.000     2.000
CH3CO              2   436.000     3.970     0.000     0.000     2.000
CH2CHO             2   436.000     3.970     0.000     0.000     2.000
CH2CO              2   436.000     3.970     0.000     0.000     2.000
HCCO               2   150.000     2.500     0.000     0.000     1.000 
CH3CO3             2   436.000     3.970     0.000     0.000     2.000
CH3CO3H            2   436.000     3.970     0.000     0.000     2.000
CH2OHCHO           2   540.215     4.796     2.730     5.200     1.000
CHOCHO             1   440.200     4.010     0.000     0.000     2.000
O2C2H4O2H          2   470.600     4.410     0.000     0.000     1.500
HO2CH2CHO          2   275.049     5.428     0.000     0.000     1.000
CH3OCHO            2   395.000     4.037     1.300     0.000     1.000
CH3OCO             2   395.000     4.037     1.300     0.000     1.000
C3H8               2   303.400     4.810     0.000     0.000     1.000
IC3H7              2   303.400     4.810     0.000     0.000     1.000
NC3H7              2   303.400     4.810     0.000     0.000     1.000
C3H6               2   307.800     4.140     0.000     0.000     1.000
C3H5-A             2   316.000     4.220     0.000     0.000     1.000
C3H5-S             2   316.000     4.220     0.000     0.000     1.000
C3H5-T             2   316.000     4.220     0.000     0.000     1.000
C3H5O              2   424.600     4.820     0.000     0.000     1.000
C3H6O              2   411.000     4.820     0.000     0.000     1.000
CH3CHCHO           2   387.860     4.687     0.000     0.000     0.000
AC4H7OOH           2   330.435     5.741     0.000     0.000     1.000
CH3CHCO            2   443.200     4.120     0.000     0.000     1.000
AC3H5OOH           2   481.500     4.997     1.700     0.000     1.000
C3H6OH1-2          2   487.900     4.820     0.000     0.000     1.000
C3H6OH2-1          2   487.900     4.820     0.000     0.000     1.000
HOC3H6O2           2   487.900     4.820     0.000     0.000     1.000
SC3H5OH            2   304.276     5.450     0.000     0.000     1.000
C3H5OH             2   481.500     4.997     1.700     0.000     1.000
CH2CCH2OH          2   481.500     4.997     1.700     0.000     1.000
C3H4-P             1   324.800     4.290     0.000     0.000     1.000
C3H4-A             1   324.800     4.290     0.000     0.000     1.000
C3H3               1   324.800     4.290     0.000     0.000     1.000
C3H2               2   209.000     4.100     0.000     0.000     1.000
C2H5CHO            2   435.200     4.662     2.700     0.000     1.000
CH2CH2CHO          2   424.600     4.820     0.000     0.000     1.000
RALD3	           2   411.000     4.820     0.000     0.000     1.000
C2H3CHO            2   443.200     4.120     0.000     0.000     1.000
CH3COCH3           2   411.000     4.820     0.000     0.000     1.000
CH3COCH2           2   424.600     4.820     0.000     0.000     1.000
NC4H10             2   352.000     5.240     0.000     0.000     1.000
PC4H9              2   352.000     5.240     0.000     0.000     1.000
SC4H9              2   352.000     5.240     0.000     0.000     1.000
IC4H10             2   335.700     5.208     0.100     0.000     1.000
IC4H9              2   352.000     5.240     0.000     0.000     1.000
TC4H9              2   352.000     5.240     0.000     0.000     1.000
IC4H8              2   344.500     5.089     0.500     0.000     1.000
IC4H7              2   355.000     4.650     0.000     0.000     1.000
IC4H7O             2   496.000     5.200     0.000     0.000     1.000
C4H8-1             2   355.000     4.650     0.000     0.000     1.000
C4H8-2             2   355.000     4.650     0.000     0.000     1.000
C4H71-3            2   357.100     4.720     0.000     0.000     1.000
C4H71-4            2   357.100     4.720     0.000     0.000     1.000
C4H71-O            2   496.000     5.200     0.000     0.000     1.000
C4H6               2   357.000     4.720     0.000     0.000     1.000
C4H5               2   357.000     5.180     0.000     0.000     1.000
C4H4               2   357.000     5.180     0.000     0.000     1.000
C4H3               1   357.000     5.180     0.000     0.000     1.000 
C4H2               1   357.000     5.180     0.000     0.000     1.000
C6H6               2   468.500     5.230     0.000     10.30     1.000
FULVENE            2   468.500     5.230     0.000     0.000     1.000
C6H5               2   412.300     5.349     0.000     0.000     1.000
C5H6               1   408.000     5.200     0.000     0.000     1.000
C5H5               1   408.000     5.200     0.000     0.000     1.000
MCPTD              2   408.000     5.200     0.000     0.000     1.000
C10H8              2   630.400     6.180     0.000     16.50     1.000
NO                 1    97.500     3.621     0.000     1.760     4.000  
N2O                1   232.400     3.828     0.000     0.000     1.000                              
NO2                2   200.000     3.500     0.000     0.000     1.000                              
HNO                2   116.700     3.492     0.000     0.000     1.000
HNO2               2   200.000     3.500     0.000     0.000     1.000                              
HONO               2   200.000     3.500     0.000     0.000     1.000                              
HONO2              2   300.000     3.500     0.000     0.000     1.000                              
N2H2               2    71.400     3.798     0.000     0.000     1.000
H2NN               2    71.400     3.798     0.000     0.000     1.000
NH2OH              2   116.700     3.492     0.000     0.000     1.000
HNOH               2   116.700     3.492     0.000     0.000     1.000
NH3                2   481.000     2.920     1.470     0.000    10.000
N2H4               2   205.000     4.230     0.000     4.260     1.500
N                  0    71.400     3.298     0.000     0.000     0.000                              
NO3                2   300.000     3.500     0.000     0.000     1.000                              
NH                 1    80.000     2.650     0.000     0.000     4.000                              
NNH                2    71.400     3.798     0.000     0.000     1.000                              
NH2                2    80.000     2.650     0.000     2.260     4.000                              
H2NO               2   116.700     3.492     0.000     0.000     1.000                              
N2H3               2   200.000     3.900     0.000     0.000     1.000
HCN                1   569.000     3.630     0.000     0.000     1.000 
HNC                1   569.000     3.630     0.000     0.000     1.000
HNCO               2   232.400     3.828     0.000     0.000     1.000 
HCNO               2   232.400     3.828     0.000     0.000     1.000                              
HOCN               2   232.400     3.828     0.000     0.000     1.000
CH2NO              2   232.400     3.828     0.000     0.000     1.000
CH3NO              1    97.500     3.621     0.000     1.760     4.000
CH3NO2             2   200.000     4.500     0.000     0.000     1.000
CH3ONO             2   200.000     4.500     0.000     0.000     1.000
CH3ONO2            2   300.000     4.500     0.000     0.000     1.000
CH3CN              1   500.000     4.630     0.000     0.000     1.000
CN                 1    75.000     3.856     0.000     0.000     1.000
NCN                1   232.400     3.828     0.000     0.000     1.000
NCO                1   232.400     3.828     0.000     0.000     1.000
HNCN		   1   232.400	   3.828     0.000     0.000     1.000
H2CN               1   569.000     3.630     0.000     0.000     1.000
HCNH               1   569.000     3.630     0.000     0.000     1.000
C2N2		   1   349.000	   4.361     0.000     0.000     1.000
CH2CN              1   232.400     3.828     0.000     0.000     1.000
CH2NH              2   417.000     3.690     1.700     0.000     2.000
CH3NH2             2   481.800     3.626     0.000     0.000     1.000
CH2NH2             2   481.800     3.626     0.000     0.000     1.000
CH3NH              2   481.800     3.626     0.000     0.000     1.000
C4H5N		   2   357.000     5.180     0.000     0.000     1.000
PYRLNE             2   357.000     5.180     0.000     0.000     1.000
PYRLYL             2   357.000     5.180     0.000     0.000     1.000
HNCPROP            2   357.000     5.180     0.000     0.000     1.000
A-C3H4CN           2   357.000     5.180     0.000     0.000     1.000
C-C3H4CN           2   357.000     5.180     0.000     0.000     1.000
C3H4CN		   2   357.000     5.180     0.000     0.000     1.000
A-C3H5CN	   2   357.000     5.180     0.000     0.000     1.000
C-C3H5CN	   2   357.000     5.180     0.000     0.000     1.000
T-C3H5CN	   2   357.000     5.180     0.000     0.000     1.000
CHCHCN             2   290.616     4.368     0.000     0.000     1.000
CH2CHCN            2   290.616     4.368     0.000     0.000     1.000
C3HN		   1   324.800     4.290     0.000     0.000     1.000
C4H4N2		   2   357.000     5.180     0.000     0.000     1.000
C4H3N2		   2   357.000     5.180     0.000     0.000     1.000
C4H2N2		   2   357.000     5.180     0.000     0.000     1.000
C2H5CN		   2   357.000     5.180     0.000     0.000     1.000
CH2CH2CN	   2   357.000     5.180     0.000     0.000     1.000
CH3CHCN 	   2   357.000     5.180     0.000     0.000     1.000
CH2N		   2   238.400     3.496     0.000     0.000     1.500
HCCN               0   311.187     4.135     0.000     0.000     0.000
C2N		   2   238.400     3.496     0.000     0.000     1.500
C4N2		   2   357.000     5.180     0.000     0.000     1.000
PYRLYLO            0   478.875     5.285     0.000     0.000     0.000
PYRLYLOOH          0   534.141     5.623     0.000     0.000     0.000
C4H4NO             0   478.875     5.285     0.000     0.000     0.000
PYRLYLOO           0   530.983     5.605     0.000     0.000     0.000
CH2CCHCN           0   418.538     4.895     0.000     0.000     0.000
C4H3NOLR           0   475.456     5.263     0.000     0.000     0.000
A-C3H4CNOOH        0   534.141     5.623     0.000     0.000     0.000
NCCO               0   375.740     4.603     0.000     0.000     0.000
OCHCN              0   379.790     4.632     0.000     0.000     0.000
OCH2CN             0   383.809     4.659     0.000     0.000     0.000
CH2NO2             0   399.427     4.766     0.000     0.000     0.000 ! FM approx
CHCNH              0   315.823     4.170     0.000     0.000     0.000 ! FM approx
C4H4N              0   422.286     4.920     0.000     0.000     0.000 ! FM approx
LC4H4N             0   422.286     4.920     0.000     0.000     0.000 ! FM approx
C4H5NOH            0   485.662     5.327     0.000     0.000     0.000 ! FM approx
C4H4NOH            0   482.278     5.306     0.000     0.000     0.000 ! FM approx
C4H3NOH            0   478.875     5.285     0.000     0.000     0.000 ! FM approx
LC4H5NOH           0   485.662     5.327     0.000     0.000     0.000 ! FM approx
AC4H4NO            0   478.875     5.285     0.000     0.000     0.000 ! FM approx
OC4H3NO            0   527.811     5.585     0.000     0.000     0.000 ! FM approx
HNC3H3CHO          0   482.278     5.306     0.000     0.000     0.000 ! FM approx
OC4H4NOH           0   534.141     5.623     0.000     0.000     0.000 ! FM approx
OC4H3NOH           0   530.983     5.605     0.000     0.000     0.000 ! FM approx
HOC4H5NO           0   537.286     5.642     0.000     0.000     0.000 ! FM approx
HOC4H5NOOH         0   588.484     5.942     0.000     0.000     0.000 ! FM approx
C4H3NO             0   475.456     5.263     0.000     0.000     0.000 ! FM approx
