! This thermodynamic database was obtained by fitting the thermodynamic properties
! extracted from the following file: CHEMKIN/Coal_NO_120.therm
! The thermodynamic properties are fitted in order to preserve not only the 
! continuity of each function at the intermediate temperature, but also the  continuity
! of the derivatives, from the 1st to the 3rd order
! The intermediate temperatures are chosen in order to minimize the fitting error.
! Last update: 11/3/2021

THERMO ALL
   270.   1000.   3500. 
N2                      N   2               G    200.00   3500.00 1050.00      1
 2.81166073e+00 1.67067353e-03-6.79997428e-07 1.32881379e-10-1.02767442e-14    2
-8.69811580e+02 6.64838050e+00 3.73100682e+00-1.83159730e-03 4.32324661e-06    3
-3.04378151e-09 7.46071562e-13-1.06287426e+03 2.16821198e+00                   4
H2                      H   2               G    200.00   3500.00  700.00      1
 3.78199881e+00-1.01873260e-03 1.24226233e-06-4.19011899e-10 4.75543794e-14    2
-1.10283023e+03-5.60525910e+00 2.64204438e+00 5.49529275e-03-1.27163634e-05    3
 1.28749174e-08-4.70027750e-12-9.43236613e+02-5.12231094e-01                   4
H                       H   1               G    200.00   3500.00  860.00      1
 2.50031493e+00-7.73406872e-07 6.39345384e-10-2.12551804e-13 2.44479207e-17    2
 2.54736474e+04-4.48357228e-01 2.49950544e+00 2.99164057e-06-5.92759783e-09    3
 4.87810185e-12-1.45539326e-15 2.54737866e+04-4.44574018e-01                   4
O2                      O   2               G    200.00   3500.00  700.00      1
 2.82012408e+00 2.48211357e-03-1.51202094e-06 4.48556202e-10-4.87305668e-14    2
-9.31350148e+02 7.94914552e+00 3.74403921e+00-2.79740148e-03 9.80122560e-06    3
-1.03259643e-08 3.79931247e-12-1.06069827e+03 3.82132645e+00                   4
O                       O   1               G    200.00   3500.00  720.00      1
 2.62549143e+00-2.08959648e-04 1.33918549e-07-3.85875908e-11 4.38918703e-15    2
 2.92061519e+04 4.48358518e+00 3.14799201e+00-3.11174063e-03 6.18137893e-06    3
-5.63808794e-09 1.94866014e-12 2.91309118e+04 2.13446550e+00                   4
H2O                     H   2O   1          G    200.00   3500.00 1420.00      1
 2.66777075e+00 3.05768849e-03-9.00442411e-07 1.43361552e-10-1.00857817e-14    2
-2.98875645e+04 6.91191131e+00 4.06061172e+00-8.65807189e-04 3.24409528e-06    3
-1.80243079e-09 3.32483293e-13-3.02831314e+04-2.96150481e-01                   4
OH                      H   1O   1          G    200.00   3500.00 1700.00      1
 2.49867369e+00 1.66635279e-03-6.28251516e-07 1.28346806e-10-1.05735894e-14    2
 3.88110716e+03 7.78218863e+00 3.91354631e+00-1.66275926e-03 2.30920029e-06    3
-1.02359508e-09 1.58829629e-13 3.40005047e+03 2.05474719e-01                   4
H2O2                    H   2O   2          G    200.00   3500.00 1800.00      1
 4.76869639e+00 3.89237848e-03-1.21382349e-06 1.92615285e-10-1.22581990e-14    2
-1.80900220e+04-5.11811777e-01 3.34774224e+00 7.05005437e-03-3.84522006e-06    3
 1.16720661e-09-1.47618105e-13-1.75784785e+04 7.17868851e+00                   4
HO2                     H   1O   2          G    200.00   3500.00  700.00      1
 3.02391889e+00 4.46390907e-03-2.23146492e-06 6.12710800e-10-6.64266237e-14    2
 3.99341609e+02 9.10699973e+00 3.61994299e+00 1.05805704e-03 5.06678942e-06    3
-6.33800762e-09 2.41597281e-12 3.15898234e+02 6.44411482e+00                   4
CO                      C   1O   1          G    200.00   3500.00  960.00      1
 2.79255381e+00 1.87486886e-03-8.59711925e-07 1.91200070e-10-1.67855286e-14    2
-1.41723335e+04 7.41443560e+00 3.75723891e+00-2.14465241e-03 5.42079004e-06    3
-4.17025963e-09 1.11901127e-12-1.43575530e+04 2.79976799e+00                   4
CO2                     C   1O   2          G    200.00   3500.00 1450.00      1
 4.70876468e+00 2.62914704e-03-9.30606462e-07 1.43892920e-10-7.62581413e-15    2
-4.90562639e+04-2.34976452e+00 2.31684347e+00 9.22755036e-03-7.75654093e-06    3
 3.28225360e-09-5.48722482e-13-4.83626067e+04 1.00786234e+01                   4
CH4                     C   1H   4          G    300.00   3500.00  700.00      1
 5.05346456e-01 1.23697844e-02-4.99807911e-06 1.04392761e-09-8.62897368e-14    2
-9.58982503e+03 1.61752773e+01 5.23967310e+00-1.46835107e-02 5.29732676e-05    3
-5.41668788e-08 1.96318554e-11-1.02526308e+04-4.97649641e+00                   4
CH3                     C   1H   3          G    300.00   3500.00 1060.00      1
 2.78805104e+00 6.15233477e-03-2.21179349e-06 3.74402648e-10-2.48151348e-14    2
 1.65862829e+04 5.77899817e+00 3.47829310e+00 3.54764774e-03 1.47408439e-06    3
-1.94375954e-09 5.21921230e-13 1.64399516e+04 2.40875956e+00                   4
CH2                     C   1H   2          G    300.00   3500.00 1800.00      1
 2.81272972e+00 3.55431388e-03-1.28768523e-06 2.21273744e-10-1.48738147e-14    2
 4.62073492e+04 6.64284652e+00 3.76489460e+00 1.43839191e-03 4.75583077e-07    3
-4.31788591e-10 7.58292874e-14 4.58645699e+04 1.48953153e+00                   4
CH2S                    C   1H   2          G    300.00   3500.00  970.00      1
 2.75934299e+00 3.65468306e-03-1.35589913e-06 2.74980408e-10-2.36795469e-14    2
 5.06429079e+04 6.11646381e+00 4.18185434e+00-2.21134312e-03 7.71527537e-06    3
-5.95950378e-09 1.58314628e-12 5.03669407e+04-7.03002582e-01                   4
CH3O                    C   1H   3O   1     G    300.00   3500.00 1740.00      1
 5.72238062e+00 5.90227638e-03-1.80340720e-06 2.13335010e-10-5.61816419e-15    2
-7.86252217e+01-7.49173676e+00 8.89660986e-01 1.70119767e-02-1.13807350e-05    3
 3.88280928e-09-5.32841479e-13 1.60316121e+03 1.85001134e+01                   4
CH2O                    C   1H   2O   1     G    300.00   3500.00  700.00      1
 1.33335655e+00 1.00905182e-02-5.12952555e-06 1.25425205e-09-1.19639106e-13    2
-1.39080170e+04 1.59916142e+01 4.32621280e+00-7.01151756e-03 3.15176939e-05    3
-3.36478617e-08 1.23454015e-11-1.43270169e+04 2.62028968e+00                   4
HCO                     C   1H   1O   1     G    200.00   3500.00  770.00      1
 2.60049318e+00 5.29278258e-03-2.69184211e-06 7.21357799e-10-7.43521409e-14    2
 4.05725330e+03 1.07450933e+01 4.03483979e+00-2.15836864e-03 1.18233875e-05    3
-1.18459406e-08 4.00593955e-12 3.83636392e+03 4.20008770e+00                   4
C2H6                    C   2H   6          G    300.00   3500.00 1800.00      1
 4.07959141e+00 1.57445262e-02-5.96197393e-06 1.06867182e-09-7.61012341e-14    2
-1.25948053e+04-1.43089411e+00-2.41778723e-01 2.53475709e-02-1.39645112e-05    3
 4.03257452e-09-4.87754387e-13-1.10391121e+04 2.19572625e+01                   4
C2H5                    C   2H   5          G    300.00   3500.00 1800.00      1
 5.19791360e+00 1.11042800e-02-3.71281686e-06 5.47665572e-10-2.89412605e-14    2
 1.17176215e+04-4.91382512e+00 6.75421802e-01 2.11542617e-02-1.20878017e-05    3
 3.64951180e-09-4.59753237e-13 1.33457186e+04 1.95628439e+01                   4
C2H4                    C   2H   4          G    300.00   3500.00 1650.00      1
 4.60402718e+00 9.50595350e-03-3.15129262e-06 4.53052075e-10-2.23949160e-14    2
 3.97229102e+03-3.77420904e+00-6.02932446e-02 2.08133970e-02-1.34307867e-05    3
 4.60638300e-09-6.51687481e-13 5.51151676e+03 2.10642172e+01                   4
C2H3                    C   2H   3          G    300.00   3500.00 1450.00      1
 4.18728376e+00 7.47581589e-03-2.58984227e-06 4.05265796e-10-2.35022722e-14    2
 3.38403785e+04 1.51958752e+00 1.23421214e+00 1.56222204e-02-1.10171572e-05    3
 4.27989337e-09-6.91541508e-13 3.46967692e+04 1.68637048e+01                   4
C2H2                    C   2H   2          G    300.00   3500.00  790.00      1
 4.37267451e+00 5.47212836e-03-2.03181547e-06 3.75019136e-10-2.77049085e-14    2
 2.58626598e+04-2.43835908e+00 7.70536982e-01 2.37107994e-02-3.66622035e-05    3
 2.95989753e-08-9.27579229e-12 2.64317975e+04 1.40907680e+01                   4
C2H                     C   2H   1          G    300.00   3500.00 1710.00      1
 3.41788257e+00 4.21328989e-03-1.58936946e-06 2.68739191e-10-1.73346358e-14    2
 6.72874491e+04 5.32512366e+00 4.60873599e+00 1.42766785e-03 8.54158643e-07    3
-6.83903344e-10 1.21940589e-13 6.68801772e+04-1.05894068e+00                   4
C2H5O                   C   2H   5O   1     G    300.00   3500.00  700.00      1
 1.68957253e+00 2.35453826e-02-1.23415274e-05 3.08911894e-09-2.98016650e-13    2
-3.10347953e+03 1.69410914e+01 3.27852951e+00 1.44656284e-02 7.11508866e-06    3
-1.54409916e-08 6.31987996e-12-3.32593351e+03 9.84203359e+00                   4
PC2H4OH                 C   2H   5O   1     G    300.00   3500.00 1470.00      1
 7.18479679e+00 1.17471700e-02-4.06239752e-06 6.31554727e-10-3.61645076e-14    2
-6.24418450e+03-9.60110090e+00 1.82077786e+00 2.63431399e-02-1.89562444e-05    3
 7.38613379e-09-1.18490244e-12-4.66716293e+03 1.83437446e+01                   4
CH3CHO                  C   2H   4O   1     G    300.00   3500.00 1800.00      1
 6.22195371e+00 1.06589270e-02-3.75190329e-06 6.00731629e-10-3.66603825e-14    2
-2.30621355e+04-8.31408576e+00 9.75916637e-01 2.23167871e-02-1.34667868e-05    3
 4.19883662e-09-5.36397186e-13-2.11735621e+04 2.00785613e+01                   4
CH2CHO                  C   2H   3O   1     G    300.00   3500.00 1340.00      1
 6.47703792e+00 7.91358605e-03-2.83605892e-06 4.62112658e-10-2.83231300e-14    2
-1.16170812e+03-8.37157284e+00 7.37868283e-01 2.50454357e-02-2.20135026e-05    3
 1.00031294e-08-1.80836357e-12 3.76389339e+02 2.09962836e+01                   4
CH2CO                   C   2H   2O   1     G    300.00   3500.00 1360.00      1
 5.69523628e+00 6.46841658e-03-2.33588415e-06 3.83408112e-10-2.36897851e-14    2
-8.05944305e+03-4.61154401e+00 2.49503978e+00 1.58807592e-02-1.27171444e-05    3
 5.47226118e-09-9.59140717e-13-7.18898960e+03 1.18115657e+01                   4
HCCO                    C   2H   1O   1     G    300.00   3500.00 1220.00      1
 5.81420512e+00 3.89116780e-03-1.41168609e-06 2.35668534e-10-1.49424973e-14    2
 1.94026782e+04-4.94089645e+00 3.33028661e+00 1.20351629e-02-1.14247949e-05    3
 5.70731267e-09-1.13618105e-12 2.00087543e+04 7.53650387e+00                   4
CH3OCO                  C   2H   3O   2     G    300.00   3500.00  730.00      1
 2.57527318e+00 2.11166692e-02-1.20149822e-05 3.14849389e-09-3.11411020e-13    2
-2.07588781e+04 1.60124236e+01 4.66126892e+00 9.68655559e-03 1.14715527e-05    3
-1.83003964e-08 7.03409935e-12-2.10634335e+04 6.60518521e+00                   4
C3H6                    C   3H   6          G    298.00   3500.00 1800.00      1
 6.31755201e+00 1.65820017e-02-6.59972302e-06 1.29512916e-09-1.03784375e-13    2
-3.79456071e+02-1.05616188e+01-8.55987190e-02 3.08112255e-02-1.84574096e-05    3
 5.68686491e-09-7.13747674e-13 1.92567819e+03 2.40935688e+01                   4
C3H5-A                  C   3H   5          G    298.00   3500.00 1600.00      1
 8.53877792e+00 1.04611885e-02-3.15379708e-06 3.85306883e-10-1.26413688e-14    2
 1.71766363e+04-2.28181758e+01-3.57888096e-01 3.27028536e-02-2.40053581e-05    3
 9.07345729e-09-1.37016487e-12 2.00235695e+04 2.42845603e+01                   4
C3H5O                   C   3H   5O   1     G    300.00   3500.00 1610.00      1
 9.11079978e+00 1.37589660e-02-5.15319199e-06 9.32421983e-10-6.74695911e-14    2
 7.77376170e+03-2.10036658e+01 9.27196847e-01 3.40908988e-02-2.40959865e-05    3
 8.77622923e-09-1.28545208e-12 1.04088818e+04 2.23747992e+01                   4
C3H3                    C   3H   3          G    300.00   3500.00  840.00      1
 5.75057760e+00 1.05635748e-02-4.84060957e-06 1.09040070e-09-9.80036150e-14    2
 4.00565408e+04-5.04125047e+00 1.75584152e+00 2.95861275e-02-3.88094537e-05    3
 2.80498008e-08-8.12163460e-12 4.07276565e+04 1.35345461e+01                   4
C2H3CHO                 C   3H   4O   1     G    300.00   3500.00 1600.00      1
 9.22597838e+00 1.12038372e-02-3.67974366e-06 5.08180254e-10-2.25803378e-14    2
-1.23719484e+04-2.08137560e+01 8.18908044e-01 3.22215131e-02-2.33838148e-05    3
 8.71820988e-09-1.30539747e-12-9.68168587e+03 2.36968522e+01                   4
C4H6                    C   4H   6          G    200.00   3500.00 1800.00      1
 9.30872521e+00 1.50139591e-02-5.06688177e-06 7.84148096e-10-4.70262839e-14    2
 8.60829987e+03-2.47389586e+01 4.65225109e-01 3.46661815e-02-2.14437338e-05    3
 6.84964885e-09-8.89456944e-13 1.17919599e+04 2.31239087e+01                   4
C4H5                    C   4H   5          G    300.00   3500.00 1800.00      1
 1.90192654e+01-1.91794385e-03 4.88814513e-06-1.91833948e-09 2.24139237e-13    2
 3.48592740e+04-7.70423351e+01-2.01742307e-01 4.07954066e-02-3.07063136e-05    3
 1.12647934e-08-1.60685144e-12 4.17788367e+04 2.69857683e+01                   4
C4H4                    C   4H   4          G    300.00   3500.00 1290.00      1
 7.65777119e+00 1.26498258e-02-4.62248952e-06 7.81217086e-10-5.07629111e-14    2
 3.13366016e+04-1.49692661e+01 7.13119719e-01 3.41836288e-02-2.96617953e-05    3
 1.37214268e-08-2.55855549e-12 3.31283217e+04 2.03030643e+01                   4
C6H6                    C   6H   6          G    300.00   3500.00 1410.00      1
 1.15055544e+01 1.99961046e-02-7.07935462e-06 1.10673029e-09-6.24178906e-14    2
 4.11452291e+03-4.24445090e+01-6.99882110e+00 7.24907868e-02-6.29247613e-05    3
 2.75111779e-08-4.74405754e-12 9.33275680e+03 5.31863191e+01                   4
FULVENE                 C   6H   6          G    200.00   3500.00 1560.00      1
 1.44152220e+01 1.47750067e-02-3.90939181e-06 2.82308156e-10 1.62511622e-14    2
 1.91167581e+04-5.54965184e+01-3.67012639e+00 6.11476948e-02-4.84985149e-05    3
 1.93374890e-08-3.03746371e-12 2.47593868e+04 3.97971310e+01                   4
C6H5                    C   6H   5          G    300.00   3500.00 1390.00      1
 1.12331261e+01 1.77269650e-02-6.33615685e-06 1.00236866e-09-5.75481757e-14    2
 3.49856300e+04-3.80075864e+01-6.76261385e+00 6.95132669e-02-6.22206553e-05    3
 2.78054854e-08-4.87825263e-12 3.99884457e+04 5.47375207e+01                   4
C5H6                    C   5H   6          G    200.00   3500.00 1630.00      1
 1.35786764e+01 1.28174257e-02-3.11961936e-06 1.29368392e-10 2.76958521e-14    2
 9.43770579e+03-5.26289052e+01-4.05866643e+00 5.60992486e-02-4.29495178e-05    3
 1.64197154e-08-2.47082363e-12 1.51874796e+04 4.10783319e+01                   4
C5H5                    C   5H   5          G    300.00   3500.00  700.00      1
 4.01652580e+00 2.68451889e-02-1.26423017e-05 2.78092329e-09-2.35299432e-13    2
 2.91110159e+04 1.44025771e+00-2.58737429e+00 6.45817609e-02-9.35063844e-05    3
 7.97943354e-08-2.77400895e-11 3.00355619e+04 3.09448125e+01                   4
MCPTD                   C   6H   8          G    300.00   3500.00 1800.00      1
-1.21144536e+02 2.92206055e-01-1.95445895e-04 5.59670227e-08-5.79656645e-12    2
 5.40571676e+04 6.85330263e+02 7.45334886e+00 6.43297727e-03 4.26983361e-05    3
-3.22345445e-08 6.45365122e-12 7.76192896e+03-1.06683176e+01                   4
C10H8                   C  10H   8          G    300.00   3500.00 1370.00      1
 1.51184828e+01 3.89675576e-02-1.78248658e-05 3.92092279e-09-3.39215689e-13    2
 1.01121562e+04-6.09041102e+01-8.71832426e+00 1.08564074e-01-9.40254318e-05    3
 4.10014902e-08-7.10574258e-12 1.66434413e+04 6.15987877e+01                   4
CYC5H4O                 C   5H   4O   1     G    300.00   3500.00 1260.00      1
 6.34459579e+00 2.39841575e-02-8.32755387e-06 8.47127652e-10 2.86249485e-14    2
 3.08659308e+03-9.73181555e+00-5.14379339e+00 6.04552343e-02-5.17455024e-05    3
 2.38195872e-08-4.52940274e-12 5.98166715e+03 4.83481227e+01                   4
C6H4O2                  C   6H   4O   2     G    300.00   3500.00 1410.00      1
 1.74929577e+01 1.29021286e-02-2.02976642e-06-3.72417846e-10 8.59745728e-14    2
-2.22100459e+04-6.49015838e+01-5.23446578e+00 7.73770890e-02-7.06201498e-05    3
 3.20580235e-08-5.66410367e-12-1.58009124e+04 5.25540058e+01                   4
CRESOL                  C   7H   8O   1     G    300.00   3500.00 1310.00      1
 1.22673687e+01 3.34155283e-02-1.38949871e-05 2.56768166e-09-1.71519559e-13    2
-2.17187243e+04-3.95715124e+01-4.41843936e+00 8.43645604e-02-7.22335735e-05    3
 3.22565297e-08-5.83733025e-12-1.73470426e+04 4.54334869e+01                   4
RCRESOLC                C   7H   7O   1     G    300.00   3500.00 1150.00      1
 1.31541709e+01 2.50657189e-02-5.32353913e-06-2.12687588e-10 1.25840459e-13    2
-3.38086418e+03-4.22339552e+01-6.42956805e+00 9.31830717e-02-9.41722601e-05    3
 5.12938173e-08-1.10712258e-11 1.12339577e+03 5.49833260e+01                   4
RCRESOLO                C   7H   7O   1     G    300.00   3500.00 1150.00      1
 1.27824815e+01 2.40796404e-02-4.51347916e-06-4.25076440e-10 1.44988501e-13    2
-3.97704756e+03-4.00543788e+01-6.60757189e+00 9.15233042e-02-9.24834755e-05    3
 5.05720229e-08-1.09413374e-11 4.82664707e+02 5.62014116e+01                   4
C6H5C2H                 C   8H   6          G    200.00   3500.00 1280.00      1
 1.52608076e+01 2.33328927e-02-9.12947229e-06 1.67060897e-09-1.19620450e-13    2
 3.14643486e+04-5.61979008e+01-2.98097334e+00 8.03384582e-02-7.59328693e-05    3
 3.64640449e-08-6.91521341e-12 3.61342445e+04 3.63113150e+01                   4
C6H4C2H                 C   8H   5          G    200.00   3500.00 1410.00      1
 1.60102852e+01 1.80276839e-02-6.10631287e-06 8.89485624e-10-4.39310920e-14    2
 6.01004863e+04-5.91795508e+01-2.59308039e+00 7.08031891e-02-6.22504674e-05    3
 2.74351852e-08-4.75061541e-12 6.53466354e+04 3.69628594e+01                   4
C6H5C2H3                C   8H   8          G    200.00   3500.00 1620.00      1
 2.08689853e+01 1.76153525e-02-4.02709967e-06 7.62333198e-11 4.96213073e-14    2
 7.92336685e+03-8.97908225e+01-4.75261288e+00 8.08785579e-02-6.26041417e-05    3
 2.41820119e-08-3.67040626e-12 1.62247647e+04 4.61791070e+01                   4
C6H5C2H2                C   8H   7          G    200.00   3500.00 1520.00      1
 1.92541493e+01 1.80154928e-02-5.00513523e-06 4.35360010e-10 9.55509219e-15    2
 3.83998804e+04-7.81182474e+01-4.29898225e+00 7.99974179e-02-6.61715087e-05    3
 2.72627168e-08-4.40283911e-12 4.55600324e+04 4.53739369e+01                   4
INDENE                  C   9H   8          G    200.00   3500.00 1610.00      1
 2.31048443e+01 1.91297591e-02-4.53548120e-06 1.22196710e-10 5.15078704e-14    2
 8.53092089e+03-1.04304478e+02-6.87762290e+00 9.36203608e-02-7.39366630e-05    3
 2.88597461e-08-4.41084452e-12 1.81852753e+04 5.46222708e+01                   4
INDENYL                 C   9H   7          G    200.00   3500.00 1430.00      1
 2.02650248e+01 2.20602643e-02-7.28401475e-06 9.93375838e-10-4.12199482e-14    2
 2.49669757e+04-8.59379552e+01-6.82385337e+00 9.78333502e-02-8.67662727e-05    3
 3.80480416e-08-6.51930836e-12 3.27143949e+04 5.44392228e+01                   4
C10H7                   C  10H   7          G    200.00   3500.00 1490.00      1
 2.12397127e+01 2.27484190e-02-6.96640085e-06 8.04033892e-10-1.68765826e-14    2
 3.76445830e+04-9.11799918e+01-6.45168838e+00 9.70877508e-02-8.18046543e-05    3
 3.42887110e-08-5.63511100e-12 4.58966205e+04 5.34576808e+01                   4
C10H7OH                 C  10H   8O   1     G    300.00   3500.00 1730.00      1
 2.61818224e+01 2.47079229e-02-8.75472975e-06 1.41213209e-09-8.61580367e-14    2
-1.58338687e+04-1.19314317e+02-3.09194614e+00 9.23929369e-02-6.74411581e-05    3
 2.40273261e-08-3.35424965e-12-5.70514482e+03 3.79602738e+01                   4
C10H7O                  C  10H   7O   1     G    200.00   3500.00 1520.00      1
 2.51245261e+01 2.12349446e-02-5.95579175e-06 5.14900720e-10 1.27936894e-14    2
 2.27944423e+03-1.11444345e+02-6.17635896e+00 1.03605695e-01-8.72427162e-05    3
 3.61670606e-08-5.85104839e-12 1.17949133e+04 5.26703358e+01                   4
C14H9                   C  14H   9          G    298.15   3500.00 1380.00      1
 2.51054797e+01 4.12375740e-02-1.71094086e-05 3.35330088e-09-2.55891933e-13    2
 4.20489547e+04-1.12231126e+02-1.15966330e+01 1.47620510e-01-1.32743034e-04    3
 5.92149558e-08-1.03757569e-11 5.21787378e+04 7.66564973e+01                   4
C16H10                  C  16H  10          G    200.00   3500.00 1560.00      1
 3.81807346e+01 2.83119223e-02-6.73305412e-06 1.57165250e-10 8.21178663e-14    2
 9.09208909e+03-1.88517714e+02-1.17161985e+01 1.56252776e-01-1.29753106e-04    3
 5.27298370e-08-8.34298979e-12 2.46599322e+04 7.43946040e+01                   4
C16H9                   C  16H   9          G    300.00   3500.00 1240.00      1
 1.61933977e+01 6.96117135e-02-3.71054121e-05 9.43826013e-09-9.32515879e-13    2
 4.61008358e+04-6.54256237e+01-1.33382684e+01 1.64875153e-01-1.52343443e-04    3
 7.13941909e-08-1.34236310e-11 5.34246890e+04 8.34001920e+01                   4
C6H5OH                  C   6H   6O   1     G    300.00   3500.00 1430.00      1
 1.28001859e+01 2.34800709e-02-9.95091013e-06 2.04936550e-09-1.68127257e-13    2
-1.75399709e+04-4.51377556e+01-4.57275686e+00 7.20757150e-02-6.09253620e-05    3
 2.58136787e-08-4.32272747e-12-1.25713093e+04 4.48905084e+01                   4
C6H5CHO                 C   7H   6O   1     G    200.00   3500.00 1630.00      1
 2.06104936e+01 1.34209230e-02-2.83635978e-06-5.48103783e-11 5.23167108e-14    2
-1.43315560e+04-8.70895599e+01-3.50845143e+00 7.26085180e-02-5.73034718e-05    3
 2.22221271e-08-3.36439149e-12-6.46877992e+03 4.10544422e+01                   4
C6H5CO                  C   7H   5O   1     G    300.00   3500.00 1470.00      1
 1.31799087e+01 2.42895707e-02-1.09067387e-05 2.35371847e-09-2.00195165e-13    2
 5.86598787e+03-4.37756649e+01-1.56203256e+00 6.44036967e-02-5.18395203e-05    3
 2.09173383e-08-3.35727336e-12 1.02001186e+04 3.30251959e+01                   4
C7H7                    C   7H   7          G    200.00   3500.00 1600.00      1
 1.77148781e+01 1.72901839e-02-4.74309316e-06 3.88421745e-10 1.27959347e-14    2
 1.68881058e+04-7.24712964e+01-3.23806381e+00 6.96725387e-02-5.38515508e-05    3
 2.08502791e-08-3.18436927e-12 2.35930472e+04 3.84624951e+01                   4
CH3C6H4                 C   7H   7          G    200.00   3500.00 1730.00      1
 1.83842182e+01 1.52647348e-02-3.43004338e-06 5.73661648e-11 4.21798063e-14    2
 2.84624024e+04-7.44700925e+01-2.82564598e+00 6.43048832e-02-4.59504033e-05    3
 1.64428613e-08-2.32566631e-12 3.58010154e+04 3.94808224e+01                   4
C6H5O                   H   5C   6O   1     G    100.00   3500.00 1800.00      1
 1.20320192e+01 2.29423311e-02-1.10171059e-05 2.53057377e-09-2.25735901e-13    2
 2.17286270e+02-4.10084348e+01 4.06305309e-01 4.87772509e-02-3.25462057e-05    3
 1.05043144e-08-1.33319988e-12 4.40254327e+03 2.19123540e+01                   4
C6H5O2                  C   6H   5O   2     G    300.00   3500.00 1300.00      1
 1.17436568e+01 2.50264983e-02-1.11158434e-05 2.39771212e-09-2.04780347e-13    2
 1.03023085e+04-3.29345583e+01-2.98072562e+00 7.03322902e-02-6.33917572e-05    3
 2.92058730e-08-5.36019591e-12 1.41306479e+04 4.19652270e+01                   4
OOC6H4OH                H   5C   6O   3     G    100.00   3500.00 1570.00      1
 2.76569225e+01 2.91346362e-04 5.46428411e-06-2.09157763e-09 2.40972769e-13    2
-1.39658759e+04-1.18517523e+02-4.81896279e-01 7.19826044e-02-6.30305484e-05    3
 2.69932769e-08-4.39037350e-12-5.13028675e+03 2.99287472e+01                   4
C6H4OH                  C   6H   5O   1     G    300.00   3500.00 1170.00      1
 1.35501563e+01 1.98692226e-02-8.43356665e-06 1.70584597e-09-1.35582640e-13    2
 1.32571078e+04-4.75538960e+01-6.19433347e+00 8.73717518e-02-9.49752707e-05    3
 5.10173582e-08-1.06722306e-11 1.78773184e+04 5.08018127e+01                   4
BZFUR                   C   8H   6O   1     G    300.00   3500.00 1380.00      1
 1.64578334e+01 2.37623566e-02-8.52218598e-06 1.36123710e-09-7.97159889e-14    2
-5.90596972e+03-6.59480381e+01-8.70136947e+00 9.66875823e-02-8.77887356e-05    3
 3.96542563e-08-7.01685714e-12 1.03797027e+03 6.35339364e+01                   4
TETRALIN                C  10H  12          G    300.00   3500.00 1650.00      1
 2.40250678e+01 3.45031690e-02-1.26565535e-05 2.20632462e-09-1.51941205e-13    2
-9.85314331e+03-1.11161770e+02-1.00807336e+01 1.17183900e-01-8.78208542e-05    3
 3.25757390e-08-4.75336763e-12 1.40177116e+03 7.04583499e+01                   4
RTETRALIN               C  10H  11          G    300.00   3500.00 1800.00      1
 2.92428061e+01 2.67835937e-02-9.17249481e-06 1.42952536e-09-8.46466182e-14    2
 3.95646504e+03-1.44540610e+02-1.09331575e+01 1.16063513e-01-8.35724273e-05    3
 2.89850559e-08-3.91180364e-12 1.84198119e+04 7.29000859e+01                   4
RTETRAOO                C  10H  11O   2     G    300.00   3500.00 1800.00      1
 5.34619195e+01-7.89286329e-03 1.09697421e-05-3.89490432e-09 4.38586901e-13    2
-1.76924222e+04-2.71823513e+02-1.36343939e+01 1.41210055e-01-1.13282690e-04    3
 4.21245150e-08-5.95299911e-12 6.46225062e+03 9.13157315e+01                   4
C10H10                  C  10H  10          G    300.00   3500.00 1800.00      1
 1.82592698e+01 4.15934216e-02-1.83631832e-05 3.88491135e-09-3.27420808e-13    2
 4.39687821e+03-8.23923218e+01-1.14588964e+01 1.07633791e-01-7.33968243e-05    3
 2.42677414e-08-3.15836943e-12 1.50954180e+04 7.84485932e+01                   4
NO                      N   1O   1          G    200.00   3500.00  800.00      1
 2.84621514e+00 2.06354046e-03-1.06904715e-06 2.65706521e-10-2.54948673e-14    2
 1.00671113e+04 8.61842850e+00 4.25026596e+00-4.95671364e-03 1.20939293e-05    3
-1.07034405e-08 3.40236358e-12 9.84246312e+03 2.15799980e+00                   4
N2O                     N   2O   1          G    200.00   3500.00 1420.00      1
 4.85543722e+00 2.58052440e-03-9.33594196e-07 1.54088463e-10-9.24862860e-15    2
 8.05595827e+03-2.39060855e+00 2.51620681e+00 9.16990584e-03-7.89420840e-06    3
 3.42198245e-09-5.84582078e-13 8.72029970e+03 9.71509320e+00                   4
NO2                     N   1O   2          G    200.00   3500.00 1800.00      1
 4.19813794e+00 3.78881378e-03-2.08226003e-06 5.53837970e-10-5.45690377e-14    2
 2.49824368e+03 3.49647574e+00 2.86592221e+00 6.74929318e-03-4.54932620e-06    3
 1.46756618e-09-1.81475734e-13 2.97784134e+03 1.07067052e+01                   4
HNO                     H   1N   1O   1     G    200.00   3500.00  700.00      1
 2.88552845e+00 3.71507602e-03-9.89194577e-07 1.60505677e-10-1.61198693e-14    2
 1.18465422e+04 9.10108586e+00 4.47186928e+00-5.34972870e-03 1.84353870e-05    3
-1.83390958e-08 6.59088065e-12 1.16244545e+04 2.01371639e+00                   4
HNO2                    H   1N   1O   2     G    200.00   3500.00  700.00      1
 1.72007297e+00 1.13464166e-02-6.67663344e-06 1.82835451e-09-1.88889111e-13    2
-6.26025905e+03 1.58192354e+01 3.09881792e+00 3.46787403e-03 1.02059578e-05    3
-1.42503038e-08 5.55348886e-12-6.45328334e+03 9.65935176e+00                   4
HONO                    H   1N   1O   2     G    200.00   3500.00 1450.00      1
 5.99816567e+00 3.29505604e-03-1.07588927e-06 1.49768833e-10-6.76019596e-15    2
-1.16909495e+04-5.24156198e+00 2.71684795e+00 1.23469670e-02-1.04399351e-05    3
 4.45507726e-09-7.49054752e-13-1.07393674e+04 1.18081173e+01                   4
NH3                     H   3N   1          G    200.00   3500.00  700.00      1
 2.51781806e+00 5.95384021e-03-2.00551774e-06 3.21049857e-10-1.88806103e-14    2
-6.46278677e+03 7.18902506e+00 4.05091142e+00-2.80669328e-03 1.67670540e-05    3
-1.75575899e-08 6.36634788e-12-6.67741985e+03 3.39551794e-01                   4
N                       N   1               G    200.00   3500.00 1800.00      1
 2.42215558e+00 1.52655402e-04-9.87414150e-08 2.32518158e-11-1.22034408e-15    2
 5.61344054e+04 4.62162566e+00 2.50554288e+00-3.26497078e-05 5.56795096e-08    3
-3.39411193e-11 6.72311912e-15 5.61043859e+04 4.17031620e+00                   4
NH                      H   1N   1          G    200.00   3500.00 1670.00      1
 2.48662839e+00 1.81565444e-03-7.12541166e-07 1.51936873e-10-1.23899449e-14    2
 4.24864648e+04 7.43461547e+00 3.66298286e+00-1.00196106e-03 1.81825120e-06    3
-8.58359483e-10 1.38852024e-13 4.20935624e+04 1.15612276e+00                   4
NH2                     N   1H   2          G    200.00   3500.00 1280.00      1
 2.55273412e+00 3.54675597e-03-1.12718085e-06 1.61534507e-10-6.97197513e-15    2
 2.15912601e+04 8.13032012e+00 4.10678625e+00-1.30965693e-03 4.56392802e-06    3
-2.80258469e-09 5.71957556e-13 2.11934228e+04 2.49283504e-01                   4
H2NO                    N   1H   2O   1     G    200.00   3500.00  700.00      1
 2.72801504e+00 7.40936630e-03-3.46220929e-06 8.08344165e-10-7.54853119e-14    2
 6.86495538e+03 9.84388852e+00 3.66110547e+00 2.07742096e-03 7.96338786e-06    3
-1.00731769e-08 3.81077222e-12 6.73432272e+03 5.67507654e+00                   4
HCN                     C   1H   1N   1     G    200.00   3500.00  780.00      1
 3.49786301e+00 3.76915269e-03-1.51027204e-06 3.01080815e-10-2.43629368e-14    2
 1.43955802e+04 3.23683733e+00 2.24572677e+00 1.01903642e-02-1.38587557e-05    3
 1.08553403e-08-3.40713842e-12 1.45909135e+04 8.96656341e+00                   4
HNC                     H   1N   1C   1     G    200.00   3500.00  700.00      1
 4.41179651e+00 2.12707775e-03-4.71968004e-07 1.02353966e-12 7.69770113e-15    2
 2.16589078e+04-1.07356914e+00 2.73172541e+00 1.17274840e-02-2.10442672e-05    3
 1.95936894e-08-6.98968297e-12 2.18941178e+04 6.43256348e+00                   4
HNCO                    H   1N   1C   1O   1G    200.00   3500.00 1050.00      1
 4.68274059e+00 5.27517046e-03-2.30255409e-06 4.91740802e-10-4.20405692e-14    2
-1.59709573e+04 2.61731790e-01 2.23902625e+00 1.45845584e-02-1.56016797e-05    3
 8.93563010e-09-2.05249040e-12-1.54577773e+04 1.21704701e+01                   4
HCNO                    H   1N   1C   1O   1G    200.00   3500.00  780.00      1
 4.79767988e+00 6.41431462e-03-3.21741495e-06 7.84733929e-10-7.49876219e-14    2
 1.84217969e+04-2.20789647e+00 6.69823287e-01 2.75828100e-02-4.39260599e-05    3
 3.55784476e-08-1.12268189e-11 1.90657425e+04 1.66810126e+01                   4
CH3NO2                  C   1H   3N   1O   2G    200.00   3500.00 1800.00      1
 5.69934620e+00 1.38065607e-02-6.43453311e-06 1.45264682e-09-1.30225206e-13    2
-1.27635731e+04-5.01015009e+00 5.58676790e-01 2.52302705e-02-1.59542913e-05    3
 4.97848318e-09-6.19924700e-13-1.09129321e+04 2.28122252e+01                   4
CN                      C   1N   1          G    200.00   3500.00  890.00      1
 2.80498942e+00 1.99013249e-03-1.04863794e-06 2.95566162e-10-3.14165335e-14    2
 5.18669927e+04 7.89927658e+00 3.76469138e+00-2.32313475e-03 6.22091360e-06    3
-5.14979079e-09 1.49817812e-12 5.16961658e+04 3.38110710e+00                   4
NCO                     C   1O   1N   1     G    200.00   3500.00 1630.00      1
 5.49723499e+00 1.70371834e-03-5.14809903e-07 5.30240356e-11-1.05670803e-16    2
 1.33777864e+04-4.53940223e+00 2.90100726e+00 8.07482934e-03-6.37779548e-06    3
 2.45097315e-09-3.67889277e-13 1.42241566e+04 9.25436079e+00                   4
H2CN                    C   1H   2N   1     G    200.00   3500.00  700.00      1
 2.09516104e+00 9.19258718e-03-4.75958105e-06 1.19375090e-09-1.16674696e-13    2
 2.77113212e+04 1.25272169e+01 3.31830755e+00 2.20317853e-03 1.02177232e-05    3
-1.30703484e-08 4.97764648e-12 2.75400807e+04 7.06250773e+00                   4
CH2NH                   C   1H   3N   1     G    200.00   3500.00  700.00      1
 5.80669263e-01 1.46544725e-02-7.73860026e-06 1.97648489e-09-1.95880938e-13    2
 9.93682813e+03 1.93649676e+01 3.61447523e+00-2.68156158e-03 2.94100442e-05    3
-3.34031765e-08 1.24397124e-11 9.51209529e+03 5.81069011e+00                   4
CATECHOL                C   6H   6O   2     G    300.00   3500.00 1150.00      1
 1.43499798e+01 2.44086034e-02-1.04210956e-05 2.01938915e-09-1.47232754e-13    2
-3.94515399e+04-4.76262860e+01-5.49815263e+00 9.34455856e-02-1.00469333e-04    3
 5.42212661e-08-1.14954669e-11-3.48864694e+04 5.09034930e+01                   4
RCATEC                  C   6H   5O   2     G    300.00   3500.00 1140.00      1
 1.40810369e+01 2.16036558e-02-9.34848722e-06 1.81734388e-09-1.31737734e-13    2
-2.57458618e+04-4.55416675e+01-4.82568617e+00 8.79430349e-02-9.66371440e-05    3
 5.28633420e-08-1.13260356e-11-2.14351289e+04 4.81496571e+01                   4
C5H5N                   C   5H   5N   1     G    200.00   3500.00 1670.00      1
 1.48267817e+01 1.16940610e-02-2.71255627e-06 6.73794651e-11 3.04919610e-14    2
 9.59020019e+03-5.88760607e+01-3.87673990e+00 5.64929151e-02-4.29510479e-05    3
 1.61306496e-08-2.37418919e-12 1.58371764e+04 4.09492269e+01                   4
C5H4N                   C   5H   4N   1     G    300.00   3500.00 1200.00      1
 4.01448127e+00 3.05044876e-02-1.70734065e-05 4.57650635e-09-4.75747804e-13    2
 3.93972028e+04 4.02774415e+00-4.61416183e+00 5.92666313e-02-5.30260861e-05    3
 2.45502172e-08-4.63693757e-12 4.14680772e+04 4.72291469e+01                   4
C5H5NO                  C   5H   5N   1O   1G    300.00   3500.00 1210.00      1
 7.35479613e+00 2.90876831e-02-1.55808757e-05 3.98078705e-09-3.94557137e-13    2
 1.37527206e+04-1.40561969e+01-4.66377757e+00 6.88185053e-02-6.48339610e-05    3
 3.11174732e-08-6.00131047e-12 1.66612154e+04 4.62174586e+01                   4
C5H4NO                  C   5H   4N   1O   1G    300.00   3500.00 1210.00      1
 7.35479613e+00 2.90876831e-02-1.55808757e-05 3.98078705e-09-3.94557137e-13    2
 1.44813106e+04-1.40561969e+01-4.66377757e+00 6.88185053e-02-6.48339610e-05    3
 3.11174732e-08-6.00131047e-12 1.73898054e+04 4.62174586e+01                   4
C5H4NO2                 C   5H   4N   1O   2G    300.00   3500.00 1210.00      1
 7.35479613e+00 2.90876831e-02-1.55808757e-05 3.98078705e-09-3.94557137e-13    2
 1.44813106e+04-1.40561969e+01-4.66377757e+00 6.88185053e-02-6.48339610e-05    3
 3.11174732e-08-6.00131047e-12 1.73898054e+04 4.62174586e+01                   4
bNC4H4CO                C   5H   4N   1O   1G    300.00   3500.00 1210.00      1
 7.35479613e+00 2.90876831e-02-1.55808757e-05 3.98078705e-09-3.94557137e-13    2
 1.44813106e+04-1.40561969e+01-4.66377757e+00 6.88185053e-02-6.48339610e-05    3
 3.11174732e-08-6.00131047e-12 1.73898054e+04 4.62174586e+01                   4
C3H3ONCO                C   4H   3N   1O   2G    300.00   3500.00 1210.00      1
 7.35479613e+00 2.90876831e-02-1.55808757e-05 3.98078705e-09-3.94557137e-13    2
 1.44813106e+04-1.40561969e+01-4.66377757e+00 6.88185053e-02-6.48339610e-05    3
 3.11174732e-08-6.00131047e-12 1.73898054e+04 4.62174586e+01                   4
C4H5N                   C   4H   5N   1     G    300.00   3500.00 1270.00      1
 9.36117079e+00 1.72757987e-02-6.11652156e-06 1.06528002e-09-7.50815127e-14    2
 8.53338244e+03-2.79960862e+01-5.32461930e+00 6.35302556e-02-6.07477700e-05    3
 2.97431007e-08-5.72032180e-12 1.22635731e+04 4.63645138e+01                   4
PYRLNE                  C   4H   5N   1          300.00   3500.00  800.00      1
-2.25123907e+00 4.24713628e-02-2.50033121e-05 6.55370520e-09-6.41454366e-13    2
 1.89830569e+04 3.46894502e+01 1.18066157e+00 2.53118596e-02 7.17075637e-06    3
-2.02580185e-08 7.73720930e-12 1.84339528e+04 1.88983199e+01                   4
PYRLYL                  C   4H   4N   1     G    300.00   3500.00 1710.00      1
 1.59928065e+01 4.27268406e-03-8.46010461e-07-4.43217665e-11 2.00499051e-14    2
 2.79279746e+04-6.47967006e+01-3.55348191e+00 4.99949961e-02-4.09533017e-05    3
 1.55920491e-08-2.26596922e-12 3.46128052e+04 3.99892962e+01                   4
CH2CHCN                 C   3H   3N   1     G    200.00   3500.00 1690.00      1
 7.83484860e+00 8.38363684e-03-2.49828670e-06 2.86570364e-10-6.79796273e-15    2
 1.86233012e+04-1.71046378e+01 1.49763743e+00 2.33829532e-02-1.58112894e-05    3
 5.53824796e-09-7.83673347e-13 2.07652786e+04 1.67940584e+01                   4
CHCHCN                  C   3H   2N   1     G    200.00   3500.00 1320.00      1
 6.85861777e+00 7.74920266e-03-2.83619309e-06 4.73014718e-10-2.98345666e-14    2
 5.05394953e+04-9.37896883e+00 1.95161727e+00 2.26189012e-02-1.97335778e-05    3
 9.00704738e-09-1.64612863e-12 5.18349435e+04 1.56568112e+01                   4
C4H4CN                  C   5H   4N   1     G    200.00   3500.00 1380.00      1
 1.19289008e+01 1.36080934e-02-4.78490623e-06 7.47955845e-10-4.27746659e-14    2
 5.55441120e+04-3.26058464e+01 1.84548244e+00 4.28353929e-02-3.65537100e-05    3
 1.60952041e-08-2.82307326e-12 5.83271355e+04 1.92885209e+01                   4
CH                      C   1H   1          G    300.00   3500.00 1590.00      1
 2.27990128e+00 2.16985238e-03-7.07637884e-07 1.23973494e-10-9.56348511e-15    2
 7.11059412e+04 8.77326061e+00 3.77264332e+00-1.58547350e-03 2.83512238e-06    3
-1.36146058e-09 2.23995331e-13 7.06312492e+04 8.79407904e-01                   4
C                       C   1               G    200.00   3500.00  700.00      1
 2.49472531e+00 3.92839476e-05-6.70014980e-08 3.71818694e-11-5.07306885e-15    2
 8.54504422e+04 4.79314254e+00 2.54495192e+00-2.47725281e-04 5.48018277e-07    3
-5.48551250e-10 2.04117331e-13 8.54434105e+04 4.56874273e+00                   4
NCN                     C   1N   2          G    200.00   3500.00 1540.00      1
 6.26178527e+00 8.14604744e-04-6.32168059e-08-5.68978567e-11 1.02757866e-14    2
 5.13388447e+04-9.55046103e+00 2.82367216e+00 9.74476868e-03-8.76142843e-06    3
 3.70856172e-09-6.01000119e-13 5.23977836e+04 8.52096412e+00                   4
HNCN                    C   1H   1N   2     G    200.00   3500.00 1460.00      1
 5.71563435e+00 3.59039536e-03-1.19666899e-06 1.72409983e-10-8.44530525e-15    2
 3.58827351e+04-4.39973155e+00 3.04255635e+00 1.09138967e-02-8.72081421e-06    3
 3.60809273e-09-5.96747146e-13 3.66632738e+04 9.50791468e+00                   4
C2N2                    C   2N   2          G    200.00   3500.00  700.00      1
 5.66789416e+00 5.81681878e-03-2.89262849e-06 6.98368845e-10-6.54524514e-14    2
 3.52445641e+04-4.84945634e+00 2.74684248e+00 2.25085427e-02-3.86606082e-05    3
 3.47631115e-08-1.22314320e-11 3.56535113e+04 8.20106354e+00                   4
CH3CN                   C   2H   3N   1     G    200.00   3500.00  700.00      1
 2.04918664e+00 1.63166629e-02-8.45703420e-06 2.11771927e-09-2.06450509e-13    2
 7.64801686e+03 1.30927474e+01 3.05185722e+00 1.05871167e-02 3.82056462e-06    3
-9.57523198e-09 3.96960351e-12 7.50764298e+03 8.61306899e+00                   4
CH2CN                   C   2H   2N   1     G    200.00   3500.00 1380.00      1
 6.11859533e+00 6.12198158e-03-2.20713413e-06 3.59045101e-10-2.17707719e-14    2
 2.86608577e+04-6.42535446e+00 2.85897544e+00 1.55701552e-02-1.24768880e-05    3
 5.32027887e-09-9.20545006e-13 2.95605128e+04 1.03502971e+01                   4
HOCN                    H   1N   1C   1O   1G    200.00   3500.00 1260.00      1
 5.08605507e+00 4.40745638e-03-1.67135017e-06 3.00184383e-10-2.12769828e-14    2
-3.69516510e+03-1.53122287e+00 2.95277827e+00 1.11797637e-02-9.73362079e-06    3
 4.56593603e-09-8.67656279e-13-3.15757934e+03 9.25362984e+00                   4
AR                000000AR  1               G    300.00   5000.00 1000.00      1
 2.50000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00    2
-7.45375000E+02 4.36600000E+00 2.50000000E+00 0.00000000E+00 0.00000000E+00    3
 0.00000000E+00 0.00000000E+00-7.45375000E+02 4.36600000E+00                   4
END
